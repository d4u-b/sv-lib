//`define VERILATOR
`define RST_TIME 19
`define CK_PER   10
