//`define VERILATOR
