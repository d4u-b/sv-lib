`ifndef __FIFO_PARA_PKG_SV__
 `define __FIFO_PARA_PKG_SV__

package fifo_para_pkg;

  localparam FF_D   = 16;
  localparam FF_W   = 32;
  localparam FF_DLY = 0;

endpackage // fifo_para_pkg

`endif
